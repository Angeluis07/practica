`timescale 1ns/1ps

module eje3_tb();

// Entradas

// Salidas

eje3 UUT(
   
);



initial begin
  $dumpfile("eje3_tb.vcd");
  $dumpvars(0, eje3_tb);

  $finish;
end

endmodule