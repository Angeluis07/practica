`timescale 1ns/1ps

module eje6_tb();

// Entradas

// Salidas

//eje4 UUT(
   
//);



initial begin
  $dumpfile("eje6_tb.vcd");
  $dumpvars(0, eje6_tb);

  $finish;
end

endmodule