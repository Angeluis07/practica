///Modulo para la operación AND
module eje1(
    input wire A,
    input wire B,
    output wire X
);
    assign X = A & B;  // Operación AND entre A y B
endmodule
