`timescale 1ns/1ps

module eje4_tb();

// Entradas

// Salidas

eje4 UUT(
   
);



initial begin
  $dumpfile("eje4_tb.vcd");
  $dumpvars(0, eje4_tb);

  $finish;
end

endmodule